module install
