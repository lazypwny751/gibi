module package
