module install

import os

import pkg.package

pub fn install_packages(pkgs []string) bool {
	if pkgs.len == 0 {
		eprintln('Error: No packages specified for installation.')
		return false
	}

	for pkg in pkgs {
		if os.is_dir(pkg) {
			println('Installing package from local path: $pkg')
		} else {
			println('Installing package from remote source: $pkg')
		}
	}

	return true
}